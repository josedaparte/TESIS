** Profile: "SCHEMATIC1-flyback"  [ D:\Usuarios\josed\Documents\facu\Facu-5\potencia\DVD_Potencia2016\Diapositivas\PSPICE_cap_5\flyback-pspicefiles\schematic1\flyback.sim ] 

** Creating circuit file "flyback.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Usuarios\josed\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3m 2.5m 
.STEP PARAM load LIST 10 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
